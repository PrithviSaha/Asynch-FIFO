`define DSIZE 		8
`define num_of_txns 	20
`define ADDR 		4
`define DEPTH 		1 << `ADDR
